module alu(
    input logic[7:0]x,
    input logic[7:0]y,
    input logic[1:0]m,
    input logic[1:0]s,
    output logic[15:0]z
);
endmodule