module arithmetic(
input logic [7:0] x,
input logic [7:0] y,
input logic [1:0] m,
output logic[15:0] z);
//
endmodule