module xor2 ( 
	input logic a,   // First input 
	input logic b,   // Second input 
	output logic y   // Output 
	); 

   assign y = a ^ b;
   
endmodule