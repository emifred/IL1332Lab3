module demux4to1_module(
    input logic[7:0]x,
    input logic[1:0]s
);
endmodule